library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_0 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_0;

-- 32 kB BRAM
architecture behavioral of B_RAM_0 is

	type ram_type is array (0 to 32768) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (		0 => x"93",
		1 => x"13",
		2 => x"93",
		3 => x"13",
		4 => x"93",
		5 => x"13",
		6 => x"93",
		7 => x"13",
		8 => x"93",
		9 => x"13",
		10 => x"93",
		11 => x"13",
		12 => x"93",
		13 => x"13",
		14 => x"93",
		15 => x"13",
		16 => x"93",
		17 => x"13",
		18 => x"93",
		19 => x"13",
		20 => x"93",
		21 => x"13",
		22 => x"93",
		23 => x"13",
		24 => x"93",
		25 => x"13",
		26 => x"93",
		27 => x"13",
		28 => x"93",
		29 => x"13",
		30 => x"93",
		31 => x"93",
		32 => x"b7",
		33 => x"93",
		34 => x"37",
		35 => x"13",
		36 => x"33",
		37 => x"b7",
		38 => x"93",
		39 => x"63",
		40 => x"93",
		41 => x"b7",
		42 => x"93",
		43 => x"37",
		44 => x"13",
		45 => x"33",
		46 => x"b7",
		47 => x"93",
		48 => x"63",
		49 => x"93",
		50 => x"93",
		51 => x"13",
		52 => x"33",
		53 => x"93",
		54 => x"63",
		55 => x"93",
		56 => x"93",
		57 => x"13",
		58 => x"33",
		59 => x"93",
		60 => x"63",
		61 => x"93",
		62 => x"93",
		63 => x"13",
		64 => x"33",
		65 => x"93",
		66 => x"63",
		67 => x"93",
		68 => x"93",
		69 => x"37",
		70 => x"33",
		71 => x"93",
		72 => x"63",
		73 => x"93",
		74 => x"b7",
		75 => x"13",
		76 => x"33",
		77 => x"93",
		78 => x"63",
		79 => x"93",
		80 => x"b7",
		81 => x"37",
		82 => x"33",
		83 => x"93",
		84 => x"63",
		85 => x"93",
		86 => x"b7",
		87 => x"93",
		88 => x"37",
		89 => x"13",
		90 => x"33",
		91 => x"b7",
		92 => x"93",
		93 => x"63",
		94 => x"93",
		95 => x"b7",
		96 => x"93",
		97 => x"37",
		98 => x"13",
		99 => x"33",
		100 => x"b7",
		101 => x"93",
		102 => x"63",
		103 => x"93",
		104 => x"b7",
		105 => x"37",
		106 => x"33",
		107 => x"93",
		108 => x"63",
		109 => x"93",
		110 => x"93",
		111 => x"13",
		112 => x"33",
		113 => x"93",
		114 => x"63",
		115 => x"93",
		116 => x"93",
		117 => x"13",
		118 => x"33",
		119 => x"93",
		120 => x"63",
		121 => x"93",
		122 => x"93",
		123 => x"13",
		124 => x"33",
		125 => x"93",
		126 => x"63",
		127 => x"93",
		128 => x"93",
		129 => x"13",
		130 => x"b3",
		131 => x"93",
		132 => x"63",
		133 => x"93",
		134 => x"93",
		135 => x"13",
		136 => x"33",
		137 => x"93",
		138 => x"63",
		139 => x"93",
		140 => x"93",
		141 => x"b3",
		142 => x"93",
		143 => x"63",
		144 => x"93",
		145 => x"13",
		146 => x"93",
		147 => x"13",
		148 => x"33",
		149 => x"13",
		150 => x"13",
		151 => x"93",
		152 => x"e3",
		153 => x"93",
		154 => x"63",
		155 => x"93",
		156 => x"13",
		157 => x"93",
		158 => x"13",
		159 => x"33",
		160 => x"13",
		161 => x"13",
		162 => x"13",
		163 => x"93",
		164 => x"e3",
		165 => x"93",
		166 => x"63",
		167 => x"93",
		168 => x"13",
		169 => x"93",
		170 => x"13",
		171 => x"33",
		172 => x"13",
		173 => x"13",
		174 => x"13",
		175 => x"13",
		176 => x"93",
		177 => x"e3",
		178 => x"93",
		179 => x"63",
		180 => x"93",
		181 => x"13",
		182 => x"93",
		183 => x"13",
		184 => x"33",
		185 => x"13",
		186 => x"93",
		187 => x"e3",
		188 => x"93",
		189 => x"63",
		190 => x"93",
		191 => x"13",
		192 => x"93",
		193 => x"13",
		194 => x"13",
		195 => x"33",
		196 => x"13",
		197 => x"93",
		198 => x"e3",
		199 => x"93",
		200 => x"63",
		201 => x"93",
		202 => x"13",
		203 => x"93",
		204 => x"13",
		205 => x"13",
		206 => x"13",
		207 => x"33",
		208 => x"13",
		209 => x"93",
		210 => x"e3",
		211 => x"93",
		212 => x"63",
		213 => x"93",
		214 => x"13",
		215 => x"93",
		216 => x"13",
		217 => x"13",
		218 => x"33",
		219 => x"13",
		220 => x"93",
		221 => x"e3",
		222 => x"93",
		223 => x"63",
		224 => x"93",
		225 => x"13",
		226 => x"93",
		227 => x"13",
		228 => x"13",
		229 => x"13",
		230 => x"33",
		231 => x"13",
		232 => x"93",
		233 => x"e3",
		234 => x"93",
		235 => x"63",
		236 => x"93",
		237 => x"13",
		238 => x"93",
		239 => x"13",
		240 => x"13",
		241 => x"13",
		242 => x"33",
		243 => x"13",
		244 => x"93",
		245 => x"e3",
		246 => x"93",
		247 => x"63",
		248 => x"93",
		249 => x"13",
		250 => x"13",
		251 => x"93",
		252 => x"33",
		253 => x"13",
		254 => x"93",
		255 => x"e3",
		256 => x"93",
		257 => x"63",
		258 => x"93",
		259 => x"13",
		260 => x"13",
		261 => x"93",
		262 => x"13",
		263 => x"33",
		264 => x"13",
		265 => x"93",
		266 => x"e3",
		267 => x"93",
		268 => x"63",
		269 => x"93",
		270 => x"13",
		271 => x"13",
		272 => x"93",
		273 => x"13",
		274 => x"13",
		275 => x"33",
		276 => x"13",
		277 => x"93",
		278 => x"e3",
		279 => x"93",
		280 => x"63",
		281 => x"93",
		282 => x"13",
		283 => x"13",
		284 => x"13",
		285 => x"93",
		286 => x"33",
		287 => x"13",
		288 => x"93",
		289 => x"e3",
		290 => x"93",
		291 => x"63",
		292 => x"93",
		293 => x"13",
		294 => x"13",
		295 => x"13",
		296 => x"93",
		297 => x"13",
		298 => x"33",
		299 => x"13",
		300 => x"93",
		301 => x"e3",
		302 => x"93",
		303 => x"63",
		304 => x"93",
		305 => x"13",
		306 => x"13",
		307 => x"13",
		308 => x"13",
		309 => x"93",
		310 => x"33",
		311 => x"13",
		312 => x"93",
		313 => x"e3",
		314 => x"93",
		315 => x"63",
		316 => x"93",
		317 => x"93",
		318 => x"33",
		319 => x"93",
		320 => x"63",
		321 => x"93",
		322 => x"93",
		323 => x"33",
		324 => x"93",
		325 => x"63",
		326 => x"93",
		327 => x"b3",
		328 => x"93",
		329 => x"63",
		330 => x"93",
		331 => x"93",
		332 => x"13",
		333 => x"33",
		334 => x"93",
		335 => x"63",
		336 => x"6f",
		337 => x"b7",
		338 => x"23",
		339 => x"6f",
		340 => x"b7",
		341 => x"93",
		342 => x"23",
		343 => x"6f",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(14 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(14 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(14 downto 0))));
		end if;
	end process;

end behavioral ; -- arch