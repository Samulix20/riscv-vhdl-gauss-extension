library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_2 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_2;

-- 32 kB BRAM
architecture behavioral of B_RAM_2 is

	type ram_type is array (0 to 32768) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (		0 => x"00",
		1 => x"00",
		2 => x"00",
		3 => x"00",
		4 => x"00",
		5 => x"00",
		6 => x"00",
		7 => x"00",
		8 => x"00",
		9 => x"00",
		10 => x"00",
		11 => x"00",
		12 => x"00",
		13 => x"00",
		14 => x"00",
		15 => x"00",
		16 => x"00",
		17 => x"00",
		18 => x"00",
		19 => x"00",
		20 => x"00",
		21 => x"00",
		22 => x"00",
		23 => x"00",
		24 => x"00",
		25 => x"00",
		26 => x"00",
		27 => x"00",
		28 => x"00",
		29 => x"00",
		30 => x"00",
		31 => x"00",
		32 => x"00",
		33 => x"00",
		34 => x"db",
		35 => x"71",
		36 => x"20",
		37 => x"00",
		38 => x"03",
		39 => x"77",
		40 => x"10",
		41 => x"00",
		42 => x"00",
		43 => x"db",
		44 => x"71",
		45 => x"20",
		46 => x"00",
		47 => x"03",
		48 => x"77",
		49 => x"20",
		50 => x"00",
		51 => x"00",
		52 => x"20",
		53 => x"00",
		54 => x"77",
		55 => x"30",
		56 => x"10",
		57 => x"10",
		58 => x"20",
		59 => x"10",
		60 => x"77",
		61 => x"40",
		62 => x"30",
		63 => x"70",
		64 => x"20",
		65 => x"50",
		66 => x"77",
		67 => x"50",
		68 => x"00",
		69 => x"ff",
		70 => x"20",
		71 => x"00",
		72 => x"77",
		73 => x"60",
		74 => x"00",
		75 => x"00",
		76 => x"20",
		77 => x"00",
		78 => x"77",
		79 => x"70",
		80 => x"00",
		81 => x"ff",
		82 => x"20",
		83 => x"00",
		84 => x"77",
		85 => x"e0",
		86 => x"aa",
		87 => x"b0",
		88 => x"03",
		89 => x"d1",
		90 => x"20",
		91 => x"01",
		92 => x"f3",
		93 => x"77",
		94 => x"f0",
		95 => x"03",
		96 => x"d0",
		97 => x"aa",
		98 => x"b1",
		99 => x"20",
		100 => x"01",
		101 => x"f3",
		102 => x"77",
		103 => x"20",
		104 => x"00",
		105 => x"00",
		106 => x"20",
		107 => x"00",
		108 => x"77",
		109 => x"30",
		110 => x"f0",
		111 => x"f0",
		112 => x"20",
		113 => x"10",
		114 => x"77",
		115 => x"40",
		116 => x"f0",
		117 => x"10",
		118 => x"20",
		119 => x"f0",
		120 => x"77",
		121 => x"50",
		122 => x"10",
		123 => x"f0",
		124 => x"20",
		125 => x"f0",
		126 => x"77",
		127 => x"80",
		128 => x"d0",
		129 => x"b0",
		130 => x"20",
		131 => x"f0",
		132 => x"70",
		133 => x"90",
		134 => x"e0",
		135 => x"b0",
		136 => x"20",
		137 => x"a0",
		138 => x"71",
		139 => x"a0",
		140 => x"d0",
		141 => x"10",
		142 => x"90",
		143 => x"70",
		144 => x"b0",
		145 => x"00",
		146 => x"d0",
		147 => x"b0",
		148 => x"20",
		149 => x"07",
		150 => x"12",
		151 => x"20",
		152 => x"52",
		153 => x"f0",
		154 => x"73",
		155 => x"c0",
		156 => x"00",
		157 => x"e0",
		158 => x"b0",
		159 => x"20",
		160 => x"00",
		161 => x"07",
		162 => x"12",
		163 => x"20",
		164 => x"52",
		165 => x"a0",
		166 => x"73",
		167 => x"d0",
		168 => x"00",
		169 => x"f0",
		170 => x"b0",
		171 => x"20",
		172 => x"00",
		173 => x"00",
		174 => x"07",
		175 => x"12",
		176 => x"20",
		177 => x"52",
		178 => x"50",
		179 => x"73",
		180 => x"e0",
		181 => x"00",
		182 => x"d0",
		183 => x"b0",
		184 => x"20",
		185 => x"12",
		186 => x"20",
		187 => x"52",
		188 => x"f0",
		189 => x"77",
		190 => x"f0",
		191 => x"00",
		192 => x"e0",
		193 => x"b0",
		194 => x"00",
		195 => x"20",
		196 => x"12",
		197 => x"20",
		198 => x"52",
		199 => x"a0",
		200 => x"77",
		201 => x"00",
		202 => x"00",
		203 => x"f0",
		204 => x"b0",
		205 => x"00",
		206 => x"00",
		207 => x"20",
		208 => x"12",
		209 => x"20",
		210 => x"52",
		211 => x"50",
		212 => x"77",
		213 => x"10",
		214 => x"00",
		215 => x"d0",
		216 => x"00",
		217 => x"b0",
		218 => x"20",
		219 => x"12",
		220 => x"20",
		221 => x"52",
		222 => x"f0",
		223 => x"77",
		224 => x"20",
		225 => x"00",
		226 => x"e0",
		227 => x"00",
		228 => x"b0",
		229 => x"00",
		230 => x"20",
		231 => x"12",
		232 => x"20",
		233 => x"52",
		234 => x"a0",
		235 => x"77",
		236 => x"30",
		237 => x"00",
		238 => x"f0",
		239 => x"00",
		240 => x"00",
		241 => x"b0",
		242 => x"20",
		243 => x"12",
		244 => x"20",
		245 => x"52",
		246 => x"50",
		247 => x"77",
		248 => x"40",
		249 => x"00",
		250 => x"b0",
		251 => x"d0",
		252 => x"20",
		253 => x"12",
		254 => x"20",
		255 => x"52",
		256 => x"f0",
		257 => x"77",
		258 => x"50",
		259 => x"00",
		260 => x"b0",
		261 => x"e0",
		262 => x"00",
		263 => x"20",
		264 => x"12",
		265 => x"20",
		266 => x"52",
		267 => x"a0",
		268 => x"77",
		269 => x"60",
		270 => x"00",
		271 => x"b0",
		272 => x"f0",
		273 => x"00",
		274 => x"00",
		275 => x"20",
		276 => x"12",
		277 => x"20",
		278 => x"52",
		279 => x"50",
		280 => x"77",
		281 => x"70",
		282 => x"00",
		283 => x"b0",
		284 => x"00",
		285 => x"d0",
		286 => x"20",
		287 => x"12",
		288 => x"20",
		289 => x"52",
		290 => x"f0",
		291 => x"77",
		292 => x"80",
		293 => x"00",
		294 => x"b0",
		295 => x"00",
		296 => x"e0",
		297 => x"00",
		298 => x"20",
		299 => x"12",
		300 => x"20",
		301 => x"52",
		302 => x"a0",
		303 => x"77",
		304 => x"90",
		305 => x"00",
		306 => x"b0",
		307 => x"00",
		308 => x"00",
		309 => x"f0",
		310 => x"20",
		311 => x"12",
		312 => x"20",
		313 => x"52",
		314 => x"50",
		315 => x"77",
		316 => x"a0",
		317 => x"f0",
		318 => x"10",
		319 => x"00",
		320 => x"71",
		321 => x"b0",
		322 => x"00",
		323 => x"00",
		324 => x"00",
		325 => x"71",
		326 => x"c0",
		327 => x"00",
		328 => x"00",
		329 => x"70",
		330 => x"d0",
		331 => x"10",
		332 => x"20",
		333 => x"20",
		334 => x"00",
		335 => x"70",
		336 => x"00",
		337 => x"09",
		338 => x"30",
		339 => x"00",
		340 => x"09",
		341 => x"00",
		342 => x"30",
		343 => x"00",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(14 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(14 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(14 downto 0))));
		end if;
	end process;

end behavioral ; -- arch