library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_1 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_1;

-- 32 kB BRAM
architecture behavioral of B_RAM_1 is

	type ram_type is array (0 to 32768) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (		0 => x"00",
		1 => x"01",
		2 => x"01",
		3 => x"02",
		4 => x"02",
		5 => x"03",
		6 => x"03",
		7 => x"04",
		8 => x"04",
		9 => x"05",
		10 => x"05",
		11 => x"06",
		12 => x"06",
		13 => x"07",
		14 => x"07",
		15 => x"08",
		16 => x"08",
		17 => x"09",
		18 => x"09",
		19 => x"0a",
		20 => x"0a",
		21 => x"0b",
		22 => x"0b",
		23 => x"0c",
		24 => x"0c",
		25 => x"0d",
		26 => x"0d",
		27 => x"0e",
		28 => x"0e",
		29 => x"0f",
		30 => x"0f",
		31 => x"01",
		32 => x"80",
		33 => x"80",
		34 => x"71",
		35 => x"01",
		36 => x"87",
		37 => x"13",
		38 => x"83",
		39 => x"14",
		40 => x"01",
		41 => x"80",
		42 => x"80",
		43 => x"71",
		44 => x"01",
		45 => x"87",
		46 => x"13",
		47 => x"83",
		48 => x"12",
		49 => x"01",
		50 => x"00",
		51 => x"01",
		52 => x"87",
		53 => x"03",
		54 => x"16",
		55 => x"01",
		56 => x"00",
		57 => x"01",
		58 => x"87",
		59 => x"03",
		60 => x"1a",
		61 => x"01",
		62 => x"00",
		63 => x"01",
		64 => x"87",
		65 => x"03",
		66 => x"1e",
		67 => x"01",
		68 => x"00",
		69 => x"81",
		70 => x"87",
		71 => x"03",
		72 => x"12",
		73 => x"01",
		74 => x"00",
		75 => x"01",
		76 => x"87",
		77 => x"03",
		78 => x"16",
		79 => x"01",
		80 => x"00",
		81 => x"81",
		82 => x"87",
		83 => x"03",
		84 => x"1a",
		85 => x"01",
		86 => x"b0",
		87 => x"80",
		88 => x"01",
		89 => x"01",
		90 => x"87",
		91 => x"03",
		92 => x"83",
		93 => x"18",
		94 => x"01",
		95 => x"00",
		96 => x"80",
		97 => x"b1",
		98 => x"01",
		99 => x"87",
		100 => x"03",
		101 => x"83",
		102 => x"16",
		103 => x"01",
		104 => x"00",
		105 => x"01",
		106 => x"87",
		107 => x"03",
		108 => x"1a",
		109 => x"01",
		110 => x"00",
		111 => x"01",
		112 => x"87",
		113 => x"03",
		114 => x"1e",
		115 => x"01",
		116 => x"00",
		117 => x"01",
		118 => x"87",
		119 => x"03",
		120 => x"12",
		121 => x"01",
		122 => x"00",
		123 => x"01",
		124 => x"87",
		125 => x"03",
		126 => x"16",
		127 => x"01",
		128 => x"00",
		129 => x"01",
		130 => x"80",
		131 => x"03",
		132 => x"9a",
		133 => x"01",
		134 => x"00",
		135 => x"01",
		136 => x"81",
		137 => x"03",
		138 => x"1e",
		139 => x"01",
		140 => x"00",
		141 => x"80",
		142 => x"03",
		143 => x"94",
		144 => x"01",
		145 => x"02",
		146 => x"00",
		147 => x"01",
		148 => x"87",
		149 => x"03",
		150 => x"02",
		151 => x"02",
		152 => x"14",
		153 => x"03",
		154 => x"1e",
		155 => x"01",
		156 => x"02",
		157 => x"00",
		158 => x"01",
		159 => x"87",
		160 => x"00",
		161 => x"03",
		162 => x"02",
		163 => x"02",
		164 => x"12",
		165 => x"03",
		166 => x"16",
		167 => x"01",
		168 => x"02",
		169 => x"00",
		170 => x"01",
		171 => x"87",
		172 => x"00",
		173 => x"00",
		174 => x"03",
		175 => x"02",
		176 => x"02",
		177 => x"10",
		178 => x"03",
		179 => x"1c",
		180 => x"01",
		181 => x"02",
		182 => x"00",
		183 => x"01",
		184 => x"87",
		185 => x"02",
		186 => x"02",
		187 => x"16",
		188 => x"03",
		189 => x"18",
		190 => x"01",
		191 => x"02",
		192 => x"00",
		193 => x"01",
		194 => x"00",
		195 => x"87",
		196 => x"02",
		197 => x"02",
		198 => x"14",
		199 => x"03",
		200 => x"12",
		201 => x"01",
		202 => x"02",
		203 => x"00",
		204 => x"01",
		205 => x"00",
		206 => x"00",
		207 => x"87",
		208 => x"02",
		209 => x"02",
		210 => x"12",
		211 => x"03",
		212 => x"1a",
		213 => x"01",
		214 => x"02",
		215 => x"00",
		216 => x"00",
		217 => x"01",
		218 => x"87",
		219 => x"02",
		220 => x"02",
		221 => x"14",
		222 => x"03",
		223 => x"14",
		224 => x"01",
		225 => x"02",
		226 => x"00",
		227 => x"00",
		228 => x"01",
		229 => x"00",
		230 => x"87",
		231 => x"02",
		232 => x"02",
		233 => x"12",
		234 => x"03",
		235 => x"1c",
		236 => x"01",
		237 => x"02",
		238 => x"00",
		239 => x"00",
		240 => x"00",
		241 => x"01",
		242 => x"87",
		243 => x"02",
		244 => x"02",
		245 => x"12",
		246 => x"03",
		247 => x"14",
		248 => x"01",
		249 => x"02",
		250 => x"01",
		251 => x"00",
		252 => x"87",
		253 => x"02",
		254 => x"02",
		255 => x"16",
		256 => x"03",
		257 => x"10",
		258 => x"01",
		259 => x"02",
		260 => x"01",
		261 => x"00",
		262 => x"00",
		263 => x"87",
		264 => x"02",
		265 => x"02",
		266 => x"14",
		267 => x"03",
		268 => x"1a",
		269 => x"01",
		270 => x"02",
		271 => x"01",
		272 => x"00",
		273 => x"00",
		274 => x"00",
		275 => x"87",
		276 => x"02",
		277 => x"02",
		278 => x"12",
		279 => x"03",
		280 => x"12",
		281 => x"01",
		282 => x"02",
		283 => x"01",
		284 => x"00",
		285 => x"00",
		286 => x"87",
		287 => x"02",
		288 => x"02",
		289 => x"14",
		290 => x"03",
		291 => x"1c",
		292 => x"01",
		293 => x"02",
		294 => x"01",
		295 => x"00",
		296 => x"00",
		297 => x"00",
		298 => x"87",
		299 => x"02",
		300 => x"02",
		301 => x"12",
		302 => x"03",
		303 => x"14",
		304 => x"01",
		305 => x"02",
		306 => x"01",
		307 => x"00",
		308 => x"00",
		309 => x"00",
		310 => x"87",
		311 => x"02",
		312 => x"02",
		313 => x"12",
		314 => x"03",
		315 => x"1c",
		316 => x"01",
		317 => x"00",
		318 => x"01",
		319 => x"03",
		320 => x"12",
		321 => x"01",
		322 => x"00",
		323 => x"81",
		324 => x"03",
		325 => x"18",
		326 => x"01",
		327 => x"00",
		328 => x"03",
		329 => x"90",
		330 => x"01",
		331 => x"00",
		332 => x"01",
		333 => x"80",
		334 => x"03",
		335 => x"14",
		336 => x"00",
		337 => x"00",
		338 => x"a0",
		339 => x"00",
		340 => x"00",
		341 => x"01",
		342 => x"a0",
		343 => x"00",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(14 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(14 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(14 downto 0))));
		end if;
	end process;

end behavioral ; -- arch