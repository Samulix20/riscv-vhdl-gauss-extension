library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_3 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_3;

-- 32 kB BRAM
architecture behavioral of B_RAM_3 is

	type ram_type is array (0 to 32768) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (		0 => x"00",
		1 => x"00",
		2 => x"00",
		3 => x"00",
		4 => x"00",
		5 => x"00",
		6 => x"00",
		7 => x"00",
		8 => x"00",
		9 => x"00",
		10 => x"00",
		11 => x"00",
		12 => x"00",
		13 => x"00",
		14 => x"00",
		15 => x"00",
		16 => x"00",
		17 => x"00",
		18 => x"00",
		19 => x"00",
		20 => x"00",
		21 => x"00",
		22 => x"00",
		23 => x"00",
		24 => x"00",
		25 => x"00",
		26 => x"00",
		27 => x"00",
		28 => x"00",
		29 => x"00",
		30 => x"00",
		31 => x"02",
		32 => x"00",
		33 => x"e0",
		34 => x"b6",
		35 => x"db",
		36 => x"02",
		37 => x"00",
		38 => x"20",
		39 => x"4a",
		40 => x"02",
		41 => x"00",
		42 => x"fc",
		43 => x"b6",
		44 => x"db",
		45 => x"02",
		46 => x"00",
		47 => x"24",
		48 => x"48",
		49 => x"00",
		50 => x"00",
		51 => x"00",
		52 => x"02",
		53 => x"00",
		54 => x"46",
		55 => x"00",
		56 => x"00",
		57 => x"00",
		58 => x"02",
		59 => x"00",
		60 => x"44",
		61 => x"00",
		62 => x"00",
		63 => x"00",
		64 => x"02",
		65 => x"01",
		66 => x"42",
		67 => x"00",
		68 => x"00",
		69 => x"ff",
		70 => x"02",
		71 => x"00",
		72 => x"42",
		73 => x"00",
		74 => x"80",
		75 => x"00",
		76 => x"02",
		77 => x"00",
		78 => x"40",
		79 => x"00",
		80 => x"80",
		81 => x"ff",
		82 => x"02",
		83 => x"00",
		84 => x"3e",
		85 => x"01",
		86 => x"aa",
		87 => x"aa",
		88 => x"00",
		89 => x"e7",
		90 => x"02",
		91 => x"00",
		92 => x"f7",
		93 => x"3c",
		94 => x"01",
		95 => x"00",
		96 => x"e7",
		97 => x"aa",
		98 => x"aa",
		99 => x"02",
		100 => x"00",
		101 => x"f7",
		102 => x"3a",
		103 => x"02",
		104 => x"ff",
		105 => x"ff",
		106 => x"02",
		107 => x"00",
		108 => x"38",
		109 => x"02",
		110 => x"ff",
		111 => x"ff",
		112 => x"02",
		113 => x"00",
		114 => x"36",
		115 => x"02",
		116 => x"ff",
		117 => x"00",
		118 => x"02",
		119 => x"ff",
		120 => x"36",
		121 => x"02",
		122 => x"00",
		123 => x"ff",
		124 => x"02",
		125 => x"ff",
		126 => x"34",
		127 => x"00",
		128 => x"00",
		129 => x"00",
		130 => x"02",
		131 => x"08",
		132 => x"32",
		133 => x"00",
		134 => x"00",
		135 => x"00",
		136 => x"02",
		137 => x"09",
		138 => x"30",
		139 => x"00",
		140 => x"00",
		141 => x"02",
		142 => x"0a",
		143 => x"30",
		144 => x"00",
		145 => x"00",
		146 => x"00",
		147 => x"00",
		148 => x"02",
		149 => x"00",
		150 => x"00",
		151 => x"00",
		152 => x"fe",
		153 => x"08",
		154 => x"2c",
		155 => x"00",
		156 => x"00",
		157 => x"00",
		158 => x"00",
		159 => x"02",
		160 => x"00",
		161 => x"00",
		162 => x"00",
		163 => x"00",
		164 => x"fe",
		165 => x"09",
		166 => x"2a",
		167 => x"00",
		168 => x"00",
		169 => x"00",
		170 => x"00",
		171 => x"02",
		172 => x"00",
		173 => x"00",
		174 => x"00",
		175 => x"00",
		176 => x"00",
		177 => x"fe",
		178 => x"0a",
		179 => x"26",
		180 => x"00",
		181 => x"00",
		182 => x"00",
		183 => x"00",
		184 => x"02",
		185 => x"00",
		186 => x"00",
		187 => x"fe",
		188 => x"08",
		189 => x"24",
		190 => x"00",
		191 => x"00",
		192 => x"00",
		193 => x"00",
		194 => x"00",
		195 => x"02",
		196 => x"00",
		197 => x"00",
		198 => x"fe",
		199 => x"09",
		200 => x"22",
		201 => x"01",
		202 => x"00",
		203 => x"00",
		204 => x"00",
		205 => x"00",
		206 => x"00",
		207 => x"02",
		208 => x"00",
		209 => x"00",
		210 => x"fe",
		211 => x"0a",
		212 => x"1e",
		213 => x"01",
		214 => x"00",
		215 => x"00",
		216 => x"00",
		217 => x"00",
		218 => x"02",
		219 => x"00",
		220 => x"00",
		221 => x"fe",
		222 => x"08",
		223 => x"1c",
		224 => x"01",
		225 => x"00",
		226 => x"00",
		227 => x"00",
		228 => x"00",
		229 => x"00",
		230 => x"02",
		231 => x"00",
		232 => x"00",
		233 => x"fe",
		234 => x"09",
		235 => x"18",
		236 => x"01",
		237 => x"00",
		238 => x"00",
		239 => x"00",
		240 => x"00",
		241 => x"00",
		242 => x"02",
		243 => x"00",
		244 => x"00",
		245 => x"fe",
		246 => x"0a",
		247 => x"16",
		248 => x"01",
		249 => x"00",
		250 => x"00",
		251 => x"00",
		252 => x"02",
		253 => x"00",
		254 => x"00",
		255 => x"fe",
		256 => x"08",
		257 => x"14",
		258 => x"01",
		259 => x"00",
		260 => x"00",
		261 => x"00",
		262 => x"00",
		263 => x"02",
		264 => x"00",
		265 => x"00",
		266 => x"fe",
		267 => x"09",
		268 => x"10",
		269 => x"01",
		270 => x"00",
		271 => x"00",
		272 => x"00",
		273 => x"00",
		274 => x"00",
		275 => x"02",
		276 => x"00",
		277 => x"00",
		278 => x"fe",
		279 => x"0a",
		280 => x"0e",
		281 => x"01",
		282 => x"00",
		283 => x"00",
		284 => x"00",
		285 => x"00",
		286 => x"02",
		287 => x"00",
		288 => x"00",
		289 => x"fe",
		290 => x"08",
		291 => x"0a",
		292 => x"01",
		293 => x"00",
		294 => x"00",
		295 => x"00",
		296 => x"00",
		297 => x"00",
		298 => x"02",
		299 => x"00",
		300 => x"00",
		301 => x"fe",
		302 => x"09",
		303 => x"08",
		304 => x"01",
		305 => x"00",
		306 => x"00",
		307 => x"00",
		308 => x"00",
		309 => x"00",
		310 => x"02",
		311 => x"00",
		312 => x"00",
		313 => x"fe",
		314 => x"0a",
		315 => x"04",
		316 => x"01",
		317 => x"01",
		318 => x"02",
		319 => x"00",
		320 => x"04",
		321 => x"01",
		322 => x"02",
		323 => x"02",
		324 => x"00",
		325 => x"02",
		326 => x"01",
		327 => x"02",
		328 => x"00",
		329 => x"02",
		330 => x"01",
		331 => x"02",
		332 => x"02",
		333 => x"02",
		334 => x"00",
		335 => x"00",
		336 => x"01",
		337 => x"00",
		338 => x"00",
		339 => x"00",
		340 => x"00",
		341 => x"00",
		342 => x"00",
		343 => x"00",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(14 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(14 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(14 downto 0))));
		end if;
	end process;

end behavioral ; -- arch